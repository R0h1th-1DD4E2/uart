`timescale 1ns / 1ps

module framer(

    );
endmodule
